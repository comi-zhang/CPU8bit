library ieee;
use ieee.std_logic_1164.all;


entity reg_out is
    port(
        ir,pc,reg_in:  in std_logic_vector(7 downto 0);  -- ����Ĵ������ݣ�8λ
        offset,alu_a,alu_b,alu_out,reg_testa1,reg_testa2:  in std_logic_vector(7 downto 0);  -- ���� ALU ���ݣ�8λ
        reg_sel:  in std_logic_vector(1 downto 0);  -- ѡ��Ĵ����źţ�4λ
        sel:      in std_logic_vector(1 downto 0);  -- ѡ���źţ�2λ
        reg_data1,reg_data2: out std_logic_vector(7 downto 0)  -- ����Ĵ������ݣ�8λ
    );
end reg_out;

architecture behave of reg_out is
begin
    process(ir, pc, reg_in, sel, reg_sel, offset, alu_a, alu_b, alu_out, reg_testa1, reg_testa2)
    variable temp: std_logic_vector(3 downto 0);
    begin
        temp := sel & reg_sel;
        case sel is
            when "00"=>
                -- ���ѡ���ź�Ϊ "00"�����������Ĵ�������
                reg_data2 <= reg_in;
            when "01"=>
                -- ���ѡ���ź�Ϊ "01"�������ѡ��ļĴ����ź������Ӧ������
                case reg_sel is
                    when "00"=>
                        reg_data2 <= offset;
                    when "01"=>
                        reg_data2 <= alu_a;
                    when "10"=>
                        reg_data2 <= alu_b;
                    when "11"=>
                        reg_data2 <= alu_out;
                end case;
            when "10"=>
				case reg_sel is
                    when "00"=>
                        reg_data2 <= pc;
                    when "01"=>
                        reg_data2 <= ir;
                    when others=>
						reg_data2 <= (others => '0');  -- ����������������ȫ��
                end case;
            when "11"=>
                -- ���ѡ���ź�Ϊ "11"�������ѡ��ļĴ����ź������Ӧ������
                case reg_sel is
                    when "00"=>
						reg_data1 <= reg_testa1;
                        reg_data2 <= reg_testa2;
                    when others=>
                        reg_data2 <= (others => '0');  -- ����������������ȫ��
                end case;
            when others=>
                reg_data2 <= (others => '0');  -- ��������ѡ���ź�ֵ�����ȫ��
        end case;
    end process;
end behave;
